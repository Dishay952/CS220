module JohnsonCounter_tb;

  JohnsonCounter 

  initial begin
    begin
      $finish;
    end
  end


endmodule
